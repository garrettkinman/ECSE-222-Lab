library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity g34_clock_divider is
	port (	enable	: in	std_logic;
				reset		: in	std_logic;
				clk		: in	std_logic;
				en_out	: out	std_logic);
end g34_clock_divider;


architecture a1 of g34_clock_divider is
	-- TODO: architecture
	-- TODO: process


end a1;